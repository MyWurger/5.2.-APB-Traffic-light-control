module svetofor
#(parameter CONTROL_REG_ADDR = 4'h0,    // адрес контрольного регистра
  parameter CURRENT_STATE_ADDR = 4'h4)  // адрес регистра текущего состояния

(
    input wire PWRITE,            // сигнал, выбирающий режим записи или чтения (1 - запись, 0 - чтение)
    input wire PCLK,              // сигнал синхронизации
    input wire PSEL,              // сигнал выбора периферии 
    input wire [31:0] PADDR,      // адрес регистра
    input wire [31:0] PWDATA,     // данные для записи в регистр
    input wire PENABLE,           // сигнал разрешения
    output reg [31:0] PRDATA = 0, // данные, прочитанные из регистра
    output reg PREADY = 0         // сигнал готовности (флаг того, что всё сделано успешно)
);


reg CONTROL_REG = 0;              // контрольный регистр изначально обнулён
reg [3:0] current_state = 0;      // регистр тукущего состояния изначально обнулён


// определим набор состояний системы для перехода в разные из них на основе временных интервалов
typedef enum logic [2:0] 
{
    STATE_0,
    STATE_1,
    STATE_2,
    STATE_3,
    STATE_4,
    STATE_5
} state_t;

// временные интервалы для каждого состояния контроллера светофора. 
// Эти параметры представляют количество тактовых циклов, которые должно длиться каждое
// состояние перед переходом в следующее состояние
 
parameter TIME_STATE_0 = 15;    // 100 тактов
parameter TIME_STATE_1 = 5;     // 10 тактов
parameter TIME_STATE_2 = 5;     // 10 тактов
parameter TIME_STATE_3 = 15;    // 100 тактов
parameter TIME_STATE_4 = 5;     // 10 тактов
parameter TIME_STATE_5 = 5;     // 10 тактов
parameter TIME_STATE_6 = 15;    // 100 тактов

// Устанавливаем начальное состояние системы светофоров как STATE_0
state_t state = STATE_0;

// Определяем переменную счетчика, которая используется для отслеживания временных интервалов
// для каждого состояния контроллера светофора
// Если счетчик достигает требуемого интервала времени, функция переходит в следующее состояние и сбрасывает счетчик в 0
logic [31:0] counter = 0;


// Эти параметры представляют собой двоичные значения, которые используются для управления
// светофорами в каждом состоянии
parameter RED = 2'b00;        // красный цвет
parameter YELLOW = 2'b01;     // жёлтый цвет
parameter GREEN = 2'b10;      // зелёный цвет


// Определение различных состояний светофора для каждого направления в контроллере светофора
logic [3:0] state_0 = {GREEN, RED};     // состояние ЗЕЛЕНОЕ для первого светофора и КРАСНОЕ для второго
logic [3:0] state_1 = {YELLOW, RED};    // состояние ЖЕЛТЫЙ для первого светофора и КРАСНЫЙ для второго
logic [3:0] state_2 = {RED, YELLOW};    // состояние КРАСНЫЙ для первого светофора и ЖЁЛТЫЙ для второго
logic [3:0] state_3 = {RED, GREEN};     // состояние КРАСНЫЙ для первого светофора и ЗЕЛЁНЫЙ для второго

// определение операции со светофором и установка контрольного регистра
// при положительном фронте сигнала PCLK
always @(posedge PCLK) 
begin
    // запрос на чтение: выбрано переферийное устройство
    // сигнал записи нулевой - операция чтения
    // устройство доступно для чтения
    if (PSEL && !PWRITE && PENABLE)
     begin
        // в зависимости от того, что мы хотим прочитать
        case(PADDR)
         // чтение контрольного регистра
         CONTROL_REG_ADDR: PRDATA <= CONTROL_REG;
         // чтение регистра текущего состояния
         CURRENT_STATE_ADDR: PRDATA <= current_state;
        endcase

        // поднимаем флаг заверешения операции
        PREADY <= 1'd1;
     end

    // запрос на запись: выбрано переферийное устройство
    // сигнал записи единица - операция записи
    // устройство доступно для записи
     else if(PSEL && PWRITE && PENABLE)
     begin
        // если адрес для записи - адрес контрольного регистра
        if(PADDR == CONTROL_REG_ADDR)
         begin
            CONTROL_REG <= PWDATA;       // записываем значение в контрольный регистр
            PREADY <= 1'd1;              // поднимаем флаг заверешения операции
        end
     end
   
   // сбрасываем PREADY после выполнения записи или чтения
   if (PREADY)
    begin
      // сброс PREADY
      PREADY <= !PREADY;
    end
  end

// по негативному фронту синхросигнала убираем значение контрольного регистра
always @(negedge PCLK) 
begin
   
   // если на положительном фронте синхросигнала значение контрольного регистра
   // было установлено в высокий уровень, то устанавливаем это значение
   // в низкий уровень
   if(CONTROL_REG)
    begin
        // устанавливаем значение контрольного регистра в низкий уровень
      CONTROL_REG<=!CONTROL_REG;
    end 
end


// функция конечного автомата светофора
function void update_state();
begin

    // в зависимости от состояния светофора
    case (state)
    // ЗК
    STATE_0: begin
    // устанавливаем текущее состояние светофора
    current_state = state_0;
        if(CONTROL_REG)           // если контрольный регистр имеет значение 1, то переходим в следующее состояние принудительно
        begin
            state = STATE_1;      // устанавливаем новое состояние светофора
            counter = 0;          // сбрасываем счётчик
        end
        
        // если нет принудительного перехода в следующее состояние через управляющий регистр
        // светофор переключится в него через промежуток времени
        else if (counter == TIME_STATE_0)
        begin
            state = STATE_1;      // устанавливаем новое состояние светофора
            counter = 0;          // сбрасываем счётчик
        end
    end

    // ЖК
    STATE_1: begin
    // устанавливаем текущее состояние светофора   
    current_state = state_1;
        if(CONTROL_REG)           // если контрольный регистр имеет значение 1, то переходим в следующее состояние принудительно
        begin 
            state = STATE_2;      // устанавливаем новое состояние светофора
            counter = 0;          // сбрасываем счётчик
        end

        // если нет принудительного перехода в следующее состояние через управляющий регистр
        // светофор переключится в него через промежуток времени
        else if (counter == TIME_STATE_1)
        begin
            state = STATE_2;      // устанавливаем новое состояние светофора
            counter = 0;          // сбрасываем счётчик
        end
    end
        
    // КЖ
    STATE_2: begin
    // устанавливаем текущее состояние светофора        
    current_state = state_2;
        if(CONTROL_REG)           // если контрольный регистр имеет значение 1, то переходим в следующее состояние принудительно
        begin
            state = STATE_3;      // устанавливаем новое состояние светофора
            counter = 0;          // сбрасываем счётчик
        end

        // если нет принудительного перехода в следующее состояние через управляющий регистр
        // светофор переключится в него через промежуток времени
        else if (counter == TIME_STATE_2)
        begin
            state = STATE_3;      // устанавливаем новое состояние светофора
            counter = 0;          // сбрасываем счётчик
        end
    end

    // КЗ
    STATE_3: begin
    // устанавливаем текущее состояние светофора    
    current_state = state_3;
        if(CONTROL_REG)           // если контрольный регистр имеет значение 1, то переходим в следующее состояние принудительно
        begin
            state = STATE_4;      // устанавливаем новое состояние светофора
            counter = 0;          // сбрасываем счётчик
        end

        // если нет принудительного перехода в следующее состояние через управляющий регистр
        // светофор переключится в него через промежуток времени
        else if (counter == TIME_STATE_3)
           begin
            state = STATE_4;      // устанавливаем новое состояние светофора
            counter = 0;          // сбрасываем счётчик
          end
    end

    // КЖ
    STATE_4: begin
    // устанавливаем текущее состояние светофора 
    current_state = state_2;
        if(CONTROL_REG)           // если контрольный регистр имеет значение 1, то переходим в следующее состояние принудительно
        begin
            state = STATE_5;      // устанавливаем новое состояние светофора
            counter = 0;          // сбрасываем счётчик
        end

        // если нет принудительного перехода в следующее состояние через управляющий регистр
        // светофор переключится в него через промежуток времени
        else if (counter == TIME_STATE_4)
        begin
            state = STATE_5;      // устанавливаем новое состояние светофора
            counter = 0;          // сбрасываем счётчик
        end
    end
    
    // ЖК
    STATE_5: begin
    // устанавливаем текущее состояние светофора
    current_state = state_1;
        if(CONTROL_REG)           // если контрольный регистр имеет значение 1, то переходим в следующее состояние принудительно. возвращаемся в начало
        begin
            state = STATE_0;      // устанавливаем новое состояние светофора
            counter = 0;          // сбрасываем счётчик
        end

        // если нет принудительного перехода в следующее состояние через управляющий регистр
        // светофор переключится в него через промежуток времени
        else if (counter == TIME_STATE_5)
        begin
            state = STATE_0;      // устанавливаем новое состояние светофора. Возвращаемся в начало
            counter = 0;          // сбрасываем счётчик
        end
    end
    endcase
end
endfunction


// функция увеличения счётчика
function void increment_counter();
begin
    // увеличиваем счётчик
    counter = counter + 1;
end
endfunction


// По счётчику или высокому уровню значения контрольного регистра
always @(posedge PCLK or posedge CONTROL_REG) 
begin
    // обновляем состояние светофора
    update_state();
    // увеличиваем счётчик
    increment_counter();
end

endmodule